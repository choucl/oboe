package Config;
  typedef 64 PhysicalRegFileSize;
endpackage
