package OboeConfig;
typedef 64 NumPhysicalRegs;
Integer kNumPhysicalRegs = valueOf(NumPhysicalRegs);
endpackage
