package OboeConfig;
typedef 64 PhysicalRegFileSize;
endpackage
