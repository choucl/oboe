package OboeConfig;

// Typedef: NumPhysicalRegs
//   Number of physical registers
typedef 64 NumPhysicalRegs;

// Constant: kNumPhysicalRegs
//   Integer value of <NumPhysicalRegs>
Integer kNumPhysicalRegs = valueOf(NumPhysicalRegs);

endpackage
