package OboeConfig;

// Typedef: NumPhysicalRegs
//   Number of physical registers.
typedef 64 NumPhysicalRegs;

// Constant: kNumPhysicalRegs
//   Integer value of <NumPhysicalRegs>.
Integer kNumPhysicalRegs = valueOf(NumPhysicalRegs);

// Typedef: NumWbPorts
//   Number of write back ports
typedef 2 NumWbPorts;

// Constant: kNumWritebackPorts
//   Integer value of <NumWritebackPorts>
Integer kNumWbPorts = valueOf(NumWbPorts);

endpackage
